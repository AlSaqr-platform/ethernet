/*

Copyright (c) 2016-2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

/*
 * Generic source synchronous DDR input
 */
module ssio_ddr_in
#(
    // target ("SIM", "GENERIC", "XILINX", "ALTERA")
    parameter TARGET = "GENERIC",
    // IODDR style ("IODDR", "IODDR2")
    // Use IODDR for Virtex-4, Virtex-5, Virtex-6, 7 Series, Ultrascale
    // Use IODDR2 for Spartan-6
    parameter IODDR_STYLE = "IODDR2",
    // Clock input style ("BUFG", "BUFR", "BUFIO", "BUFIO2")
    // Use BUFR for Virtex-5, Virtex-6, 7-series
    // Use BUFG for Ultrascale
    // Use BUFIO2 for Spartan-6
    parameter CLOCK_INPUT_STYLE = "BUFIO2",
    // Width of register in bits
    parameter WIDTH = 1
)
(
    input  wire             input_clk,

    input  wire [WIDTH-1:0] input_d,

    output wire             output_clk,

    output wire [WIDTH-1:0] output_q1,
    output wire [WIDTH-1:0] output_q2
);

wire clk_int;
wire clk_io;


`ifndef GENESYSII
    generate

    if (TARGET == "XILINX") begin

        // use Xilinx clocking primitives

        if (CLOCK_INPUT_STYLE == "IBUF") begin

            // buffer RX clock

            IBUF #(
                .IBUF_LOW_PWR ("FALSE")
            )
            clk_bufio (
                .I(input_clk),
                .O(clk_int)
            );

            // pass through RX clock to logic and input buffers
            assign clk_io = clk_int;
            assign output_clk = clk_int;

        end else if (CLOCK_INPUT_STYLE == "BUFR") begin

            assign clk_int = input_clk;

            // pass through RX clock to input buffers
            BUFIO
            clk_bufio (
                .I(clk_int),
                .O(clk_io)
            );

            // pass through RX clock to logic
            BUFR #(
                .BUFR_DIVIDE("BYPASS")
            )
            clk_bufr (
                .I(clk_int),
                .O(output_clk),
                .CE(1'b1),
                .CLR(1'b0)
            );

        end else if (CLOCK_INPUT_STYLE == "BUFIO") begin

            assign clk_int = input_clk;

            // pass through RX clock to input buffers
            BUFIO
            clk_bufio (
                .I(clk_int),
                .O(clk_io)
            );

            // pass through RX clock to MAC
            BUFG
            clk_bufg (
                .I(clk_int),
                .O(output_clk)
            );

        end else if (CLOCK_INPUT_STYLE == "BUFIO2") begin

            // pass through RX clock to input buffers
            BUFIO2 #(
                .DIVIDE(1),
                .DIVIDE_BYPASS("TRUE"),
                .I_INVERT("FALSE"),
                .USE_DOUBLER("FALSE")
            )
            clk_bufio (
                .I(input_clk),
                .DIVCLK(clk_int),
                .IOCLK(clk_io),
                .SERDESSTROBE()
            );

            // pass through RX clock to MAC
            BUFG
            clk_bufg (
                .I(clk_int),
                .O(output_clk)
            );

        end

    end else begin

        // pass through RX clock to input buffers
        assign clk_io = input_clk;

        // pass through RX clock to logic
        assign clk_int = input_clk;
        assign output_clk = clk_int;

    end

    endgenerate

`else /* `ifndef GENESYSII */

    // pass through RX clock to input buffers
    assign clk_io = input_clk;

    // pass through RX clock to logic
    assign clk_int = input_clk;
    assign output_clk = clk_int;

`endif

iddr #(
    .TARGET(TARGET),
    .IODDR_STYLE(IODDR_STYLE),
    .WIDTH(WIDTH)
)
data_iddr_inst (
    .clk(clk_io),
    .d(input_d),
    .q1(output_q1),
    .q2(output_q2)
);

endmodule
