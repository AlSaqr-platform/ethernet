/*

Copyright (c) 2014-2018 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

based on fpga.v
 
*/

// Language: Verilog 2001

/*
 * RGMII top-level module
 */

module rgmii_soc (
    // Internal 125 MHz clock
    input              clk_int,
    input              rst_int,
    input              clk90_int,
    input              clk_200_int,

    /*
     * Ethernet: 1000BASE-T RGMII
     */
    input wire         phy_rx_clk,
    input wire [3:0]   phy_rxd,
    input wire         phy_rx_ctl,
    output wire        phy_tx_clk,
    output wire [3:0]  phy_txd,
    output wire        phy_tx_ctl,
    output wire        phy_reset_n,
    input wire         phy_int_n,
    input wire         phy_pme_n,
    output wire        mac_gmii_tx_en,

       /*
        * AXI input
        */
    input wire         tx_axis_tvalid,
    input wire         tx_axis_tlast,
    input wire [7:0]   tx_axis_tdata,
    output wire        tx_axis_tready,
    input wire         tx_axis_tuser,
   
       /*
        * AXI output
        */
    output wire [7:0]  rx_axis_tdata,
    output wire        rx_axis_tvalid,
    output wire        rx_axis_tlast,
    output             rx_axis_tuser,

    /*
     * Status
     */

    output wire [31:0] rx_fcs_reg,
    output wire [31:0] tx_fcs_reg

);

// IODELAY elements for RGMII interface to PHY
wire [3:0] phy_rxd_delay;
wire       phy_rx_ctl_delay;

`ifdef GENESYSII
    IDELAYCTRL idelayctrl_inst
    (
        .REFCLK(clk_200_int),
        .RST(rst_int),
        .RDY()
    );

    IDELAYE2 #(
        .IDELAY_TYPE("FIXED")
    )
    phy_rxd_idelay_0
    (
        .IDATAIN(phy_rxd[0]),
        .DATAOUT(phy_rxd_delay[0]),
        .DATAIN(1'b0),
        .C(1'b0),
        .CE(1'b0),
        .INC(1'b0),
        .CINVCTRL(1'b0),
        .CNTVALUEIN(5'd0),
        .CNTVALUEOUT(),
        .LD(1'b0),
        .LDPIPEEN(1'b0),
        .REGRST(1'b0)
    );

    IDELAYE2 #(
        .IDELAY_TYPE("FIXED")
    )
    phy_rxd_idelay_1
    (
        .IDATAIN(phy_rxd[1]),
        .DATAOUT(phy_rxd_delay[1]),
        .DATAIN(1'b0),
        .C(1'b0),
        .CE(1'b0),
        .INC(1'b0),
        .CINVCTRL(1'b0),
        .CNTVALUEIN(5'd0),
        .CNTVALUEOUT(),
        .LD(1'b0),
        .LDPIPEEN(1'b0),
        .REGRST(1'b0)
    );

    IDELAYE2 #(
        .IDELAY_TYPE("FIXED")
    )
    phy_rxd_idelay_2
    (
        .IDATAIN(phy_rxd[2]),
        .DATAOUT(phy_rxd_delay[2]),
        .DATAIN(1'b0),
        .C(1'b0),
        .CE(1'b0),
        .INC(1'b0),
        .CINVCTRL(1'b0),
        .CNTVALUEIN(5'd0),
        .CNTVALUEOUT(),
        .LD(1'b0),
        .LDPIPEEN(1'b0),
        .REGRST(1'b0)
    );

    IDELAYE2 #(
        .IDELAY_TYPE("FIXED")
    )
    phy_rxd_idelay_3
    (
        .IDATAIN(phy_rxd[3]),
        .DATAOUT(phy_rxd_delay[3]),
        .DATAIN(1'b0),
        .C(1'b0),
        .CE(1'b0),
        .INC(1'b0),
        .CINVCTRL(1'b0),
        .CNTVALUEIN(5'd0),
        .CNTVALUEOUT(),
        .LD(1'b0),
        .LDPIPEEN(1'b0),
        .REGRST(1'b0)
    );

    IDELAYE2 #(
        .IDELAY_VALUE(0),
        .IDELAY_TYPE("FIXED")
    )
    phy_rx_ctl_idelay
    (
        .IDATAIN(phy_rx_ctl),
        .DATAOUT(phy_rx_ctl_delay),
        .DATAIN(1'b0),
        .C(1'b0),
        .CE(1'b0),
        .INC(1'b0),
        .CINVCTRL(1'b0),
        .CNTVALUEIN(5'd0),
        .CNTVALUEOUT(),
        .LD(1'b0),
        .LDPIPEEN(1'b0),
        .REGRST(1'b0)
    );
`elsif FPGA_EMUL

    IDELAYCTRL #(
        .SIM_DEVICE("ULTRASCALE")
    )
    idelayctrl_inst
    (
        .REFCLK(clk_200_int),
        .RST(rst_int),
        .RDY()
    );

    generate
        genvar k;
        for(k = 0; k < 4; k++) begin
            IDELAYE3 #(
                .CASCADE("NONE"),
                .DELAY_TYPE("FIXED"),
                .REFCLK_FREQUENCY(200.0),
                .SIM_DEVICE("ULTRASCALE_PLUS")
            )
            phy_rxd_idelay_k
            (
                .CASC_OUT(),
                .CASC_IN(),
                .CASC_RETURN(),
                .IDATAIN(phy_rxd[k]),        
                .DATAOUT(phy_rxd_delay[k]),
                .DATAIN(1'b0),
                .CLK(1'b0),
                .CE(1'b0),
                .INC(1'b0),
                .CNTVALUEIN(5'd0),
                .CNTVALUEOUT(),
                .LOAD(1'b0),
                .EN_VTC(1'b1),
                .RST(1'b0)
            );
        end
    endgenerate

    /*
    IDELAYE3 #(
        .CASCADE("NONE"),
        .DELAY_TYPE("FIXED"),
        .REFCLK_FREQUENCY(200.0),
        .SIM_DEVICE("ULTRASCALE_PLUS")
    )
    phy_rxd_idelay_0
    (
        .CASC_OUT(),
        .CASC_IN(),
        .CASC_RETURN(),
        .IDATAIN(phy_rxd_ibuf[0]),        
        .DATAOUT(phy_rxd_delay[0]),
        .DATAIN(1'b0),
        .CLK(1'b0),
        .CE(1'b0),
        .INC(1'b0),
        .CNTVALUEIN(5'd0),
        .CNTVALUEOUT(),
        .LOAD(1'b0),
        .EN_VTC(1'b0),
        .RST(1'b0)
    );
    
    IDELAYE3 #(
        .CASCADE("NONE"),
        .DELAY_TYPE("FIXED"),
        .REFCLK_FREQUENCY(200.0),
        .SIM_DEVICE("ULTRASCALE_PLUS")
    )
    phy_rxd_idelay_1
    (
        .CASC_OUT(),
        .CASC_IN(),
        .CASC_RETURN(),
        .IDATAIN(phy_rxd_ibuf[1]),        
        .DATAOUT(phy_rxd_delay[1]),
        .DATAIN(1'b0),
        .CLK(1'b0),
        .CE(1'b0),
        .INC(1'b0),
        .CNTVALUEIN(5'd0),
        .CNTVALUEOUT(),
        .LOAD(1'b0),
        .EN_VTC(1'b0),
        .RST(1'b0)
    );

    IDELAYE3 #(
        .CASCADE("NONE"),
        .DELAY_TYPE("FIXED"),
        .REFCLK_FREQUENCY(200.0),
        .SIM_DEVICE("ULTRASCALE_PLUS")
    )
    phy_rxd_idelay_2
    (
        .CASC_OUT(),
        .CASC_IN(),
        .CASC_RETURN(),
        .IDATAIN(phy_rxd_ibuf[2]),        
        .DATAOUT(phy_rxd_delay[2]),
        .DATAIN(1'b0),
        .CLK(1'b0),
        .CE(1'b0),
        .INC(1'b0),
        .CNTVALUEIN(5'd0),
        .CNTVALUEOUT(),
        .LOAD(1'b0),
        .EN_VTC(1'b0),
        .RST(1'b0)
    );
    
    IDELAYE3 #(
        .CASCADE("NONE"),
        .DELAY_TYPE("FIXED"),
        .REFCLK_FREQUENCY(200.0),
        .SIM_DEVICE("ULTRASCALE_PLUS")
    )
    phy_rxd_idelay_3
    (
        .CASC_OUT(),
        .CASC_IN(),
        .CASC_RETURN(),
        .IDATAIN(phy_rxd_ibuf[3]),        
        .DATAOUT(phy_rxd_delay[3]),
        .DATAIN(1'b0),
        .CLK(1'b0),
        .CE(1'b0),
        .INC(1'b0),
        .CNTVALUEIN(5'd0),
        .CNTVALUEOUT(),
        .LOAD(1'b0),
        .EN_VTC(1'b0),
        .RST(1'b0)
    );
    */

    IDELAYE3 #(
        .CASCADE("NONE"),
        .DELAY_TYPE("FIXED"),
        .REFCLK_FREQUENCY(200.0),
        .DELAY_VALUE(0),
        .SIM_DEVICE("ULTRASCALE_PLUS")
    )
    phy_rx_ctl_idelay
    (
        .CASC_OUT(),
        .CASC_IN(),
        .CASC_RETURN(),
        .IDATAIN(phy_rx_ctl_ibuf),        
        .DATAOUT(phy_rx_ctl_delay),
        .DATAIN(1'b0),
        .CLK(1'b0),
        .CE(1'b0),
        .INC(1'b0),
        .CNTVALUEIN(5'd0),
        .CNTVALUEOUT(),
        .LOAD(1'b0),
        .EN_VTC(1'b1),
        .RST(1'b0)
    );
`else // !`ifdef GENESYSII || FPGA_EMUL
   assign phy_rx_ctl_delay = phy_rx_ctl;
   assign phy_rxd_delay = phy_rxd;
`endif

rgmii_core
core_inst (
    /*
     * Clock: 125MHz
     * Synchronous reset
     */
    .clk(clk_int),
    .clk90(clk90_int),
    .rst(rst_int),
    /*
     * Ethernet: 1000BASE-T RGMII
     */
    .phy_rx_clk(phy_rx_clk),
    .phy_rxd(phy_rxd_delay),
    .phy_rx_ctl(phy_rx_ctl_delay),
    .phy_tx_clk(phy_tx_clk),
    .phy_txd(phy_txd),
    .phy_tx_ctl(phy_tx_ctl),
    .phy_reset_n(phy_reset_n),
    .phy_int_n(phy_int_n),
    .phy_pme_n(phy_pme_n),
    .mac_gmii_tx_en(mac_gmii_tx_en),
    .tx_axis_tdata(tx_axis_tdata),
    .tx_axis_tvalid(tx_axis_tvalid),
    .tx_axis_tready(tx_axis_tready),
    .tx_axis_tlast(tx_axis_tlast),
    .tx_axis_tuser(tx_axis_tuser),
    .rx_axis_tdata(rx_axis_tdata),
    .rx_axis_tvalid(rx_axis_tvalid),
    .rx_axis_tlast(rx_axis_tlast),
    .rx_axis_tuser(rx_axis_tuser),
    .rx_fcs_reg(rx_fcs_reg),
    .tx_fcs_reg(tx_fcs_reg)
);

endmodule
